library verilog;
use verilog.vl_types.all;
entity \Multiplication__pipe_tb\ is
end \Multiplication__pipe_tb\;
