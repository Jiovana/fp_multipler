library verilog;
use verilog.vl_types.all;
entity tb_lzc8 is
end tb_lzc8;
