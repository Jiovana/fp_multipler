library verilog;
use verilog.vl_types.all;
entity Multiplication_pipe_tb is
end Multiplication_pipe_tb;
