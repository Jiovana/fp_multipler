library verilog;
use verilog.vl_types.all;
entity dequantizer_block_tb is
end dequantizer_block_tb;
