library verilog;
use verilog.vl_types.all;
entity dequantizer_block_pipe_tb is
end dequantizer_block_pipe_tb;
