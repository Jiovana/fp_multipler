library verilog;
use verilog.vl_types.all;
entity tb_int_to_fp32 is
end tb_int_to_fp32;
