library verilog;
use verilog.vl_types.all;
entity multiplication_tb_python is
end multiplication_tb_python;
