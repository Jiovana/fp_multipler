library verilog;
use verilog.vl_types.all;
entity tb_int_to_fp32_pipeline is
end tb_int_to_fp32_pipeline;
