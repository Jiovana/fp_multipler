library verilog;
use verilog.vl_types.all;
entity tb_lzc_miao_32 is
end tb_lzc_miao_32;
